library ieee;
use ieee.std_logic_1164.all;

entity ha_tb is
end ha_tb;